module Or_32(result,input1,input2);
input [31:0] input1,input2;
output [31:0] result;

or or0(result[0],input1[0],input2[0]);
or or1(result[1],input1[1],input2[1]);
or or2(result[2],input1[2],input2[2]);
or or3(result[3],input1[3],input2[3]);
or or4(result[4],input1[4],input2[4]);
or or5(result[5],input1[5],input2[5]);
or or6(result[6],input1[6],input2[6]);
or or7(result[7],input1[7],input2[7]);
or or8(result[8],input1[8],input2[8]);
or or9(result[9],input1[9],input2[9]);
or or10(result[10],input1[10],input2[10]);
or or11(result[11],input1[11],input2[11]);
or or12(result[12],input1[12],input2[12]);
or or13(result[13],input1[13],input2[13]);
or or14(result[14],input1[14],input2[14]);
or or15(result[15],input1[15],input2[15]);
or or16(result[16],input1[16],input2[16]);
or or17(result[17],input1[17],input2[17]);
or or18(result[18],input1[18],input2[18]);
or or19(result[19],input1[19],input2[19]);
or or20(result[20],input1[20],input2[20]);
or or21(result[21],input1[21],input2[21]);
or or22(result[22],input1[22],input2[22]);
or or23(result[23],input1[23],input2[23]);
or or24(result[24],input1[24],input2[24]);
or or25(result[25],input1[25],input2[25]);
or or26(result[26],input1[26],input2[26]);
or or27(result[27],input1[27],input2[27]);
or or28(result[28],input1[28],input2[28]);
or or29(result[29],input1[29],input2[29]);
or or30(result[30],input1[30],input2[30]);
or or31(result[31],input1[31],input2[31]);

endmodule